* SPICE3 file created from cmos_inv2 _3.ext - technology: scmos
.include ./t14y_tsmc_025_level3.txt
.option scale=0.1u
M1000 Vout Vin Vdd Vdd pfet w=10 l=2
+  ad=44 pd=30 as=44 ps=30
M1001 Vout Vin Gnd Gnd nfet w=5 l=2
+  ad=24 pd=20 as=24 ps=20
C0 Vdd Vin 3.3fF
C1 Gnd gnd! 12.6fF
C2 Vout gnd! 3.2fF
C3 Vin gnd! 7.7fF

vdd Vdd 0 3.3
v1 Vin 0 pulse(0 3.3 0 0.05n 0.05n 0.5n 1n)
.tran 0.01n 8n
.control
run
plot Vin Vout
.endc
end
