magic
tech scmos
timestamp 1633443764
<< nwell >>
rect -15 14 16 52
<< polysilicon >>
rect -6 41 -4 43
rect 4 41 6 43
rect -6 -10 -4 21
rect 4 -10 6 21
rect -6 -17 -4 -15
rect 4 -17 6 -15
<< ndiffusion >>
rect -8 -15 -6 -10
rect -4 -15 -2 -10
rect 2 -15 4 -10
rect 6 -15 8 -10
<< pdiffusion >>
rect -8 33 -6 41
rect -12 21 -6 33
rect -4 21 4 41
rect 6 29 12 41
rect 6 23 8 29
rect 6 21 12 23
<< metal1 >>
rect -15 50 16 52
rect -15 46 -14 50
rect -10 46 -2 50
rect 2 46 9 50
rect 13 46 16 50
rect -15 44 16 46
rect -12 41 -9 44
rect 9 19 12 23
rect -1 16 12 19
rect -1 -10 2 16
rect -12 -18 -9 -15
rect 9 -18 12 -15
rect -16 -20 15 -18
rect -16 -24 -14 -20
rect -10 -24 -4 -20
rect 0 -24 6 -20
rect 10 -24 15 -20
rect -16 -26 15 -24
<< ntransistor >>
rect -6 -15 -4 -10
rect 4 -15 6 -10
<< ptransistor >>
rect -6 21 -4 41
rect 4 21 6 41
<< polycontact >>
rect -10 4 -6 8
rect 6 3 10 7
<< ndcontact >>
rect -12 -15 -8 -10
rect -2 -15 2 -10
rect 8 -15 12 -10
<< pdcontact >>
rect -12 33 -8 41
rect 8 23 12 29
<< psubstratepcontact >>
rect -14 -24 -10 -20
rect -4 -24 0 -20
rect 6 -24 10 -20
<< nsubstratencontact >>
rect -14 46 -10 50
rect -2 46 2 50
rect 9 46 13 50
<< labels >>
rlabel polycontact -8 6 -8 6 1 X
rlabel polycontact 8 5 8 5 1 Y
rlabel metal1 -8 -23 -8 -23 1 Gnd
rlabel metal1 -6 48 -6 48 5 Vdd
rlabel metal1 11 17 11 17 1 Z
<< end >>
