magic
tech scmos
timestamp 1638005104
<< nwell >>
rect 8 70 41 71
rect 8 33 62 70
<< polysilicon >>
rect 15 58 17 60
rect 31 58 33 60
rect 15 15 17 38
rect 31 25 33 38
rect 49 27 51 29
rect 32 21 33 25
rect 31 15 33 21
rect 49 11 51 21
rect 15 3 17 5
rect 31 3 33 5
<< ndiffusion >>
rect 43 26 49 27
rect 47 22 49 26
rect 43 21 49 22
rect 51 26 57 27
rect 51 22 53 26
rect 51 21 57 22
rect 11 10 15 15
rect 14 6 15 10
rect 11 5 15 6
rect 17 10 21 15
rect 27 10 31 15
rect 17 6 18 10
rect 30 6 31 10
rect 17 5 21 6
rect 27 5 31 6
rect 33 10 37 15
rect 33 6 34 10
rect 33 5 37 6
<< pdiffusion >>
rect 11 50 15 58
rect 14 46 15 50
rect 11 38 15 46
rect 17 50 21 58
rect 27 50 31 58
rect 17 46 18 50
rect 30 46 31 50
rect 17 38 21 46
rect 27 38 31 46
rect 33 50 37 58
rect 33 46 34 50
rect 33 38 37 46
<< metal1 >>
rect 8 68 62 71
rect 8 64 19 68
rect 23 64 31 68
rect 35 64 62 68
rect 8 63 62 64
rect 10 50 13 63
rect 26 50 29 63
rect 19 25 22 46
rect 35 25 38 46
rect 19 22 28 25
rect 19 10 22 22
rect 35 22 43 25
rect 35 10 38 22
rect 10 1 13 6
rect 26 1 29 6
rect 8 0 63 1
rect 8 -4 19 0
rect 23 -4 31 0
rect 35 -4 63 0
rect 8 -7 63 -4
<< ntransistor >>
rect 49 21 51 27
rect 15 5 17 15
rect 31 5 33 15
<< ptransistor >>
rect 15 38 17 58
rect 31 38 33 58
<< polycontact >>
rect 11 21 15 25
rect 28 21 32 25
rect 51 12 55 16
<< ndcontact >>
rect 43 22 47 26
rect 53 22 57 26
rect 10 6 14 10
rect 18 6 22 10
rect 26 6 30 10
rect 34 6 38 10
<< pdcontact >>
rect 10 46 14 50
rect 18 46 22 50
rect 26 46 30 50
rect 34 46 38 50
<< psubstratepcontact >>
rect 19 -4 23 0
rect 31 -4 35 0
<< nsubstratencontact >>
rect 19 64 23 68
rect 31 64 35 68
<< psubstratepdiff >>
rect 15 -4 19 0
<< nsubstratendiff >>
rect 15 64 19 68
<< labels >>
rlabel polycontact 13 23 13 23 1 Vin
rlabel metal1 11 -2 11 -2 1 Gnd
rlabel metal1 11 66 11 66 5 Vdd
rlabel ndcontact 55 24 55 24 7 Vout
rlabel polycontact 53 14 53 14 7 clock
<< end >>
