magic
tech scmos
timestamp 1633491284
<< nwell >>
rect -40 40 38 78
<< polysilicon >>
rect -31 70 -29 72
rect -21 70 -19 72
rect -11 70 -9 72
rect 17 60 19 62
rect -31 16 -29 40
rect -21 16 -19 40
rect -11 16 -9 40
rect 17 17 19 50
rect -31 9 -29 11
rect -21 9 -19 11
rect -11 9 -9 11
rect 17 10 19 12
<< ndiffusion >>
rect -33 11 -31 16
rect -29 11 -27 16
rect -23 11 -21 16
rect -19 11 -17 16
rect -13 11 -11 16
rect -9 11 -7 16
rect 16 13 17 17
rect 13 12 17 13
rect 19 13 20 17
rect 19 12 23 13
<< pdiffusion >>
rect -39 63 -31 70
rect -34 57 -31 63
rect -39 40 -31 57
rect -29 40 -21 70
rect -19 40 -11 70
rect -9 51 -3 70
rect 13 57 17 60
rect 16 53 17 57
rect -9 45 -7 51
rect 13 50 17 53
rect 19 57 23 60
rect 19 53 20 57
rect 19 50 23 53
rect -9 40 -3 45
<< metal1 >>
rect -40 74 -39 78
rect -35 74 -27 78
rect -23 74 -17 78
rect -13 74 -7 78
rect -3 75 38 78
rect -3 74 5 75
rect -40 71 5 74
rect 9 71 17 75
rect 21 71 28 75
rect 32 71 38 75
rect -40 70 38 71
rect -40 63 -37 70
rect 12 57 15 70
rect -6 31 -3 45
rect -6 28 13 31
rect -6 24 -3 28
rect -27 21 -3 24
rect -27 16 -24 21
rect -6 16 -3 21
rect 21 17 24 53
rect -37 8 -34 11
rect -16 8 -13 11
rect 12 8 15 13
rect -38 7 38 8
rect -34 3 -26 7
rect -22 3 -15 7
rect -11 3 -4 7
rect 0 3 5 7
rect 9 3 17 7
rect 21 3 27 7
rect 31 3 38 7
rect -38 0 38 3
<< ntransistor >>
rect -31 11 -29 16
rect -21 11 -19 16
rect -11 11 -9 16
rect 17 12 19 17
<< ptransistor >>
rect -31 40 -29 70
rect -21 40 -19 70
rect -11 40 -9 70
rect 17 50 19 60
<< polycontact >>
rect -36 27 -31 32
rect -26 27 -21 32
rect -16 27 -11 32
rect 13 28 17 32
<< ndcontact >>
rect -37 11 -33 16
rect -27 11 -23 16
rect -17 11 -13 16
rect -7 11 -3 16
rect 12 13 16 17
rect 20 13 24 17
<< pdcontact >>
rect -40 57 -34 63
rect 12 53 16 57
rect -7 45 -1 51
rect 20 53 24 57
<< psubstratepcontact >>
rect -38 3 -34 7
rect -26 3 -22 7
rect -15 3 -11 7
rect -4 3 0 7
rect 5 3 9 7
rect 17 3 21 7
rect 27 3 31 7
<< nsubstratencontact >>
rect -39 74 -35 78
rect -27 74 -23 78
rect -17 74 -13 78
rect -7 74 -3 78
rect 5 71 9 75
rect 17 71 21 75
rect 28 71 32 75
<< labels >>
rlabel metal1 13 73 13 73 5 Vdd
rlabel metal1 13 5 13 5 1 Gnd
rlabel polycontact 15 30 15 30 1 Vin
rlabel polycontact -34 29 -34 29 3 x
rlabel polycontact -24 29 -24 29 1 y
rlabel polycontact -14 29 -14 29 1 z
rlabel metal1 23 30 23 30 1 Vout
<< end >>
