magic
tech scmos
timestamp 1633432454
<< nwell >>
rect -5 22 35 60
<< polysilicon >>
rect 5 49 7 51
rect 14 49 16 51
rect 25 49 27 51
rect 5 15 7 39
rect 14 15 16 39
rect 25 15 27 39
rect 5 -2 7 0
rect 14 -2 16 0
rect 25 -2 27 0
<< ndiffusion >>
rect -1 5 5 15
rect 3 0 5 5
rect 7 0 14 15
rect 16 0 25 15
rect 27 10 29 15
rect 27 0 33 10
<< pdiffusion >>
rect 3 44 5 49
rect -1 39 5 44
rect 7 44 14 49
rect 7 39 8 44
rect 12 39 14 44
rect 16 44 18 49
rect 22 44 25 49
rect 16 39 25 44
rect 27 44 33 49
rect 27 39 29 44
<< metal1 >>
rect -5 59 35 60
rect -5 55 -1 59
rect 3 55 8 59
rect 12 55 17 59
rect 21 55 27 59
rect 31 55 35 59
rect -5 52 35 55
rect -1 49 2 52
rect 18 49 21 52
rect 9 36 12 39
rect 9 33 22 36
rect 19 32 22 33
rect 30 32 33 39
rect 19 29 33 32
rect 30 15 33 29
rect -1 -10 2 0
rect -5 -13 35 -10
rect -5 -17 -3 -13
rect 1 -17 6 -13
rect 10 -17 17 -13
rect 21 -17 28 -13
rect 32 -17 35 -13
rect -5 -18 35 -17
<< ntransistor >>
rect 5 0 7 15
rect 14 0 16 15
rect 25 0 27 15
<< ptransistor >>
rect 5 39 7 49
rect 14 39 16 49
rect 25 39 27 49
<< polycontact >>
rect 1 30 5 34
rect 10 23 14 27
rect 21 17 25 21
<< ndcontact >>
rect -1 0 3 5
rect 29 10 33 15
<< pdcontact >>
rect -1 44 3 49
rect 8 39 12 44
rect 18 44 22 49
rect 29 39 33 44
<< psubstratepcontact >>
rect -3 -17 1 -13
rect 6 -17 10 -13
rect 17 -17 21 -13
rect 28 -17 32 -13
<< nsubstratencontact >>
rect -1 55 3 59
rect 8 55 12 59
rect 17 55 21 59
rect 27 55 31 59
<< labels >>
rlabel polycontact 23 19 23 19 1 Z
rlabel metal1 13 -15 13 -15 1 Gnd
rlabel polycontact 3 32 3 32 1 X
rlabel polycontact 12 25 12 25 1 Y
rlabel metal1 15 57 15 57 5 Vdd
rlabel metal1 31 30 31 30 7 Vout
<< end >>
