magic
tech scmos
timestamp 1633428776
<< nwell >>
rect -10 33 28 71
<< polysilicon >>
rect 7 53 9 55
rect 7 10 9 43
rect 7 3 9 5
<< ndiffusion >>
rect 6 6 7 10
rect 3 5 7 6
rect 9 6 10 10
rect 9 5 13 6
<< pdiffusion >>
rect 3 50 7 53
rect 6 46 7 50
rect 3 43 7 46
rect 9 50 13 53
rect 9 46 10 50
rect 9 43 13 46
<< metal1 >>
rect -10 68 28 71
rect -10 64 -5 68
rect -1 64 7 68
rect 11 64 18 68
rect 22 64 28 68
rect -10 63 28 64
rect 2 50 5 63
rect 11 10 14 46
rect 2 1 5 6
rect -10 0 28 1
rect -10 -4 -5 0
rect -1 -4 7 0
rect 11 -4 17 0
rect 21 -4 28 0
rect -10 -7 28 -4
<< ntransistor >>
rect 7 5 9 10
<< ptransistor >>
rect 7 43 9 53
<< polycontact >>
rect 3 21 7 25
<< ndcontact >>
rect 2 6 6 10
rect 10 6 14 10
<< pdcontact >>
rect 2 46 6 50
rect 10 46 14 50
<< psubstratepcontact >>
rect -5 -4 -1 0
rect 7 -4 11 0
rect 17 -4 21 0
<< nsubstratencontact >>
rect -5 64 -1 68
rect 7 64 11 68
rect 18 64 22 68
<< labels >>
rlabel metal1 3 66 3 66 5 Vdd
rlabel metal1 3 -2 3 -2 1 Gnd
rlabel polycontact 5 23 5 23 1 Vin
rlabel metal1 13 22 13 22 1 Vout
<< end >>
