* SPICE3 file created from cmos_nand2.ext - technology: scmos
.include ./t14y_tsmc_025_level3.txt
.option scale=0.1u

M1000 Vout X Vdd Vdd pfet w=10 l=2
+  ad=80 pd=36 as=100 ps=60
M1001 Vdd Y Vout Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_9_n18# X Gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=50 ps=30
M1003 Vout Y a_9_n18# Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 Vdd X 3.3fF
C1 Vdd Y 3.3fF
C2 Gnd gnd 9.8fF
C3 Vout gnd 3.0fF
C4 Y gnd 5.6fF
C5 X gnd 5.6fF
C7 Vout Gnd 0.1fF

vdd Vdd 0 3.3
v2 X 0 pulse(0 3.3 0 0.01n 0.01n 1n 2n)
v3 Y 0 pulse(0 3.3 0 0.01n 0.01n 2n 4n)
.tran 0.01n 4n
.control
 foreach cap 1fF 2fF 10fF 50fF 100fF 200fF 1000fF  
  alter C7=$cap 
  tran 0.01n 4n
  meas TRAN max_vout MAX V(vout)
  meas TRAN avg_power integ I(vdd) from=3n to=4n 
  PRINT avg_power*3.3/(1n)
 end
.endc

.control
let x1=-tran1.vdd#branch
let x2=-tran2.vdd#branch
let x3=-tran3.vdd#branch
let x4=-tran4.vdd#branch
let x5=-tran5.vdd#branch
let x6=-tran6.vdd#branch
let x7=-tran7.vdd#branch

let y1=tran1.Vout
let y2=tran2.Vout
let y3=tran3.Vout
let y4=tran4.Vout
let y5=tran5.Vout
let y6=tran6.Vout
let y7=tran7.Vout

plot x1 x2 x3 x4 x5 x6 x7
plot y1 y2 y3 y4 y5 y6 y7 
.endc
.end
