magic
tech scmos
timestamp 1633433652
<< nwell >>
rect 0 14 65 52
<< polysilicon >>
rect 8 34 10 36
rect 18 34 20 36
rect 44 34 46 36
rect 8 0 10 24
rect 18 0 20 24
rect 44 -9 46 24
rect 8 -12 10 -10
rect 18 -12 20 -10
rect 44 -16 46 -14
<< ndiffusion >>
rect 3 -5 8 0
rect 7 -10 8 -5
rect 10 -10 18 0
rect 20 -5 21 0
rect 20 -10 25 -5
rect 43 -13 44 -9
rect 40 -14 44 -13
rect 46 -13 47 -9
rect 46 -14 50 -13
<< pdiffusion >>
rect 7 29 8 34
rect 3 24 8 29
rect 10 29 18 34
rect 10 24 12 29
rect 16 24 18 29
rect 20 29 21 34
rect 40 31 44 34
rect 20 24 25 29
rect 43 27 44 31
rect 40 24 44 27
rect 46 31 50 34
rect 46 27 47 31
rect 46 24 50 27
<< metal1 >>
rect 0 49 65 52
rect 0 48 32 49
rect 0 44 5 48
rect 9 44 19 48
rect 23 45 32 48
rect 36 45 44 49
rect 48 45 55 49
rect 59 45 65 49
rect 23 44 65 45
rect 3 34 6 44
rect 22 34 25 44
rect 39 31 42 44
rect 13 11 16 24
rect 13 8 25 11
rect 22 6 25 8
rect 22 3 40 6
rect 22 0 25 3
rect 48 -9 51 27
rect 3 -18 6 -10
rect 39 -18 42 -13
rect 0 -19 65 -18
rect 0 -23 6 -19
rect 10 -23 18 -19
rect 22 -23 32 -19
rect 36 -23 44 -19
rect 48 -23 54 -19
rect 58 -23 65 -19
rect 0 -26 65 -23
<< ntransistor >>
rect 8 -10 10 0
rect 18 -10 20 0
rect 44 -14 46 -9
<< ptransistor >>
rect 8 24 10 34
rect 18 24 20 34
rect 44 24 46 34
<< polycontact >>
rect 4 7 8 11
rect 14 1 18 5
rect 40 2 44 6
<< ndcontact >>
rect 3 -10 7 -5
rect 21 -5 25 0
rect 39 -13 43 -9
rect 47 -13 51 -9
<< pdcontact >>
rect 3 29 7 34
rect 12 24 16 29
rect 21 29 25 34
rect 39 27 43 31
rect 47 27 51 31
<< psubstratepcontact >>
rect 6 -23 10 -19
rect 18 -23 22 -19
rect 32 -23 36 -19
rect 44 -23 48 -19
rect 54 -23 58 -19
<< nsubstratencontact >>
rect 5 44 9 48
rect 19 44 23 48
rect 32 45 36 49
rect 44 45 48 49
rect 55 45 59 49
<< labels >>
rlabel polycontact 6 9 6 9 3 X
rlabel polycontact 16 3 16 3 1 Y
rlabel metal1 12 -21 12 -21 1 Gnd
rlabel metal1 14 46 14 46 5 Vdd
rlabel metal1 50 3 50 3 1 Vout
<< end >>
