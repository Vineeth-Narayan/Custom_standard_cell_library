magic
tech scmos
timestamp 1633491915
<< nwell >>
rect -8 10 32 48
<< polysilicon >>
rect 1 40 3 42
rect 11 40 13 42
rect 21 40 23 42
rect 1 -14 3 10
rect 11 -14 13 10
rect 21 -14 23 10
rect 1 -21 3 -19
rect 11 -21 13 -19
rect 21 -21 23 -19
<< ndiffusion >>
rect -1 -19 1 -14
rect 3 -19 5 -14
rect 9 -19 11 -14
rect 13 -19 15 -14
rect 19 -19 21 -14
rect 23 -19 25 -14
<< pdiffusion >>
rect -7 33 1 40
rect -2 27 1 33
rect -7 10 1 27
rect 3 10 11 40
rect 13 10 21 40
rect 23 21 29 40
rect 23 15 25 21
rect 23 10 29 15
<< metal1 >>
rect -8 44 -7 48
rect -3 44 5 48
rect 9 44 15 48
rect 19 44 25 48
rect 29 44 30 48
rect -8 40 30 44
rect -8 33 -5 40
rect 26 -6 29 15
rect 5 -9 29 -6
rect 5 -14 8 -9
rect 26 -14 29 -9
rect -5 -22 -2 -19
rect 16 -22 19 -19
rect -6 -23 32 -22
rect -2 -27 6 -23
rect 10 -27 17 -23
rect 21 -27 28 -23
rect -6 -30 32 -27
<< ntransistor >>
rect 1 -19 3 -14
rect 11 -19 13 -14
rect 21 -19 23 -14
<< ptransistor >>
rect 1 10 3 40
rect 11 10 13 40
rect 21 10 23 40
<< polycontact >>
rect -4 -3 1 2
rect 6 -3 11 2
rect 16 -3 21 2
<< ndcontact >>
rect -5 -19 -1 -14
rect 5 -19 9 -14
rect 15 -19 19 -14
rect 25 -19 29 -14
<< pdcontact >>
rect -8 27 -2 33
rect 25 15 31 21
<< psubstratepcontact >>
rect -6 -27 -2 -23
rect 6 -27 10 -23
rect 17 -27 21 -23
rect 28 -27 32 -23
<< nsubstratencontact >>
rect -7 44 -3 48
rect 5 44 9 48
rect 15 44 19 48
rect 25 44 29 48
<< labels >>
rlabel metal1 12 46 12 46 5 Vdd
rlabel polycontact -2 -1 -2 -1 3 x
rlabel polycontact 8 -1 8 -1 1 y
rlabel polycontact 18 -1 18 -1 1 z
rlabel metal1 28 -5 28 -5 7 Vout
rlabel metal1 13 -25 13 -25 1 Gnd
<< end >>
