magic
tech scmos
timestamp 1633432035
<< nwell >>
rect -1 6 26 44
<< polysilicon >>
rect 7 26 9 28
rect 17 26 19 28
rect 7 -8 9 16
rect 17 -8 19 16
rect 7 -20 9 -18
rect 17 -20 19 -18
<< ndiffusion >>
rect 2 -13 7 -8
rect 6 -18 7 -13
rect 9 -18 17 -8
rect 19 -13 20 -8
rect 19 -18 24 -13
<< pdiffusion >>
rect 6 21 7 26
rect 2 16 7 21
rect 9 21 17 26
rect 9 16 11 21
rect 15 16 17 21
rect 19 21 20 26
rect 19 16 24 21
<< metal1 >>
rect -1 40 26 44
rect -1 36 4 40
rect 8 36 18 40
rect 22 36 26 40
rect 2 26 5 36
rect 21 26 24 36
rect 12 3 15 16
rect 12 0 24 3
rect 21 -8 24 0
rect 2 -26 5 -18
rect -1 -27 26 -26
rect -1 -31 5 -27
rect 9 -31 17 -27
rect 21 -31 26 -27
rect -1 -34 26 -31
<< ntransistor >>
rect 7 -18 9 -8
rect 17 -18 19 -8
<< ptransistor >>
rect 7 16 9 26
rect 17 16 19 26
<< polycontact >>
rect 3 -1 7 3
rect 13 -7 17 -3
<< ndcontact >>
rect 2 -18 6 -13
rect 20 -13 24 -8
<< pdcontact >>
rect 2 21 6 26
rect 11 16 15 21
rect 20 21 24 26
<< psubstratepcontact >>
rect 5 -31 9 -27
rect 17 -31 21 -27
<< nsubstratencontact >>
rect 4 36 8 40
rect 18 36 22 40
<< labels >>
rlabel polycontact 5 1 5 1 3 X
rlabel polycontact 15 -5 15 -5 1 Y
rlabel metal1 22 1 22 1 7 Vout
rlabel metal1 11 -29 11 -29 1 Gnd
rlabel metal1 13 38 13 38 5 Vdd
<< end >>
